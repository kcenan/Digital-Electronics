magic
tech scmos
timestamp 1494793225
<< nwell >>
rect -127 170 118 262
<< polysilicon >>
rect -14 257 6 275
rect -14 198 6 209
rect -14 -208 6 -178
rect -14 -237 6 -224
<< ndiffusion >>
rect -48 -212 -14 -208
rect -48 -220 -44 -212
rect -18 -220 -14 -212
rect -48 -224 -14 -220
rect 6 -212 40 -208
rect 6 -220 10 -212
rect 36 -220 40 -212
rect 6 -224 40 -220
<< pdiffusion >>
rect -48 252 -14 257
rect -48 216 -44 252
rect -21 216 -14 252
rect -48 209 -14 216
rect 6 252 40 257
rect 6 216 13 252
rect 36 216 40 252
rect 6 209 40 216
<< metal1 >>
rect -157 556 148 576
rect -118 252 -66 556
rect 58 252 110 556
rect -66 216 -44 252
rect 13 170 36 216
rect -14 47 6 170
rect 14 47 36 170
rect -92 27 6 47
rect -14 -156 6 27
rect 10 27 84 47
rect 10 -212 36 27
rect -44 -428 -18 -220
rect -44 -444 -40 -428
rect -157 -458 -40 -444
rect -22 -444 -18 -428
rect 52 -428 78 -424
rect 52 -444 56 -428
rect -22 -458 56 -444
rect 74 -444 78 -428
rect 74 -458 148 -444
rect -157 -464 148 -458
<< ntransistor >>
rect -14 -224 6 -208
<< ptransistor >>
rect -14 209 6 257
<< polycontact >>
rect -14 170 6 198
rect -14 -178 6 -156
<< ndcontact >>
rect -44 -220 -18 -212
rect 10 -220 36 -212
<< pdcontact >>
rect -44 216 -21 252
rect 13 216 36 252
<< psubstratepcontact >>
rect -40 -458 -22 -428
rect 56 -458 74 -428
<< nsubstratencontact >>
rect -118 179 -66 252
rect 58 179 110 252
<< labels >>
rlabel metal1 74 37 74 37 1 out
rlabel metal1 -88 37 -88 37 1 in
rlabel metal1 -5 566 -5 566 1 vdd!
rlabel metal1 -4 -454 -4 -454 1 gnd!
<< end >>
