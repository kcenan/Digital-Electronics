magic
tech scmos
timestamp 1494878802
<< nwell >>
rect -127 106 364 518
<< polysilicon >>
rect -14 497 6 514
rect -14 106 6 113
rect 222 497 242 504
rect 222 400 242 407
rect -14 -160 6 -152
rect -14 -299 6 -288
rect 222 -292 242 -282
rect 222 -327 242 -322
<< ndiffusion >>
rect -48 -170 -14 -160
rect -48 -280 -44 -170
rect -18 -280 -14 -170
rect -48 -288 -14 -280
rect 6 -170 40 -160
rect 6 -280 10 -170
rect 36 -280 40 -170
rect 6 -288 40 -280
rect 132 -296 222 -292
rect 132 -318 140 -296
rect 214 -318 222 -296
rect 132 -322 222 -318
rect 242 -296 330 -292
rect 242 -318 250 -296
rect 324 -318 330 -296
rect 242 -322 330 -318
<< pdiffusion >>
rect -48 474 -14 497
rect -48 120 -44 474
rect -21 120 -14 474
rect -48 113 -14 120
rect 6 474 40 497
rect 6 120 13 474
rect 36 120 40 474
rect 6 113 40 120
rect 132 486 222 497
rect 132 416 140 486
rect 214 416 222 486
rect 132 407 222 416
rect 242 486 330 497
rect 242 416 250 486
rect 324 416 330 486
rect 242 407 330 416
<< metal1 >>
rect -157 556 402 576
rect -118 502 -66 556
rect 58 502 110 556
rect 222 518 242 526
rect -66 120 -44 474
rect 13 106 36 120
rect -14 47 6 79
rect 14 47 36 106
rect -92 27 6 47
rect -92 -2 -80 16
rect -14 -28 6 27
rect -14 -128 6 -46
rect 10 27 66 47
rect 10 -170 36 27
rect 140 16 214 416
rect 140 -2 158 16
rect 184 -2 214 16
rect -44 -352 -18 -280
rect 106 -327 122 -46
rect 140 -296 214 -2
rect 250 16 324 416
rect 250 -2 364 16
rect 250 -296 324 -2
rect 106 -344 222 -327
rect -44 -357 198 -352
rect -44 -422 -31 -357
rect 189 -422 198 -357
rect -44 -428 198 -422
rect -44 -444 -40 -428
rect -157 -458 -40 -444
rect -22 -458 56 -428
rect 74 -444 198 -428
rect 74 -458 402 -444
rect -157 -464 402 -458
<< metal2 >>
rect 66 526 222 542
rect 66 47 84 526
rect -66 -2 158 16
rect 6 -46 106 -28
<< ntransistor >>
rect -14 -288 6 -160
rect 222 -322 242 -292
<< ptransistor >>
rect -14 113 6 497
rect 222 407 242 497
<< polycontact >>
rect 222 504 242 518
rect -14 79 6 106
rect -14 -152 6 -128
rect 222 -344 242 -327
<< ndcontact >>
rect -44 -280 -18 -170
rect 10 -280 36 -170
rect 140 -318 214 -296
rect 250 -318 324 -296
<< pdcontact >>
rect -44 120 -21 474
rect 13 120 36 474
rect 140 416 214 486
rect 250 416 324 486
<< m2contact >>
rect 222 526 242 542
rect -80 -2 -66 16
rect -14 -46 6 -28
rect 66 27 84 47
rect 158 -2 184 16
rect 106 -46 122 -28
<< psubstratepcontact >>
rect -31 -422 189 -357
rect -40 -458 -22 -428
rect 56 -458 74 -428
<< nsubstratencontact >>
rect -118 112 -66 502
rect 58 112 110 502
<< labels >>
rlabel metal1 -5 566 -5 566 1 vdd!
rlabel metal1 -4 -454 -4 -454 1 gnd!
rlabel metal1 -88 37 -88 37 1 S
rlabel metal1 -87 7 -87 7 1 in
rlabel metal1 359 7 359 7 1 out
<< end >>
