magic
tech scmos
timestamp 1494861522
<< nwell >>
rect -127 106 118 518
rect 373 106 618 518
rect 806 454 973 540
rect 1011 454 1170 540
<< polysilicon >>
rect 870 518 886 534
rect 930 518 946 534
rect 1038 522 1054 534
rect 1098 522 1114 534
rect -14 497 6 514
rect -14 106 6 113
rect 486 497 506 514
rect 486 106 506 113
rect 870 452 886 464
rect 930 452 946 464
rect 1038 452 1054 468
rect 1098 452 1114 468
rect -14 -160 6 -152
rect 486 -160 506 -152
rect 870 -240 886 -234
rect 930 -240 946 -234
rect 1038 -240 1054 -230
rect 1098 -240 1114 -230
rect 870 -269 886 -258
rect 930 -269 946 -258
rect 1038 -269 1054 -258
rect 1098 -269 1114 -258
rect -14 -299 6 -288
rect 486 -299 506 -288
<< ndiffusion >>
rect -48 -170 -14 -160
rect -48 -280 -44 -170
rect -18 -280 -14 -170
rect -48 -288 -14 -280
rect 6 -170 40 -160
rect 6 -280 10 -170
rect 36 -280 40 -170
rect 6 -288 40 -280
rect 452 -170 486 -160
rect 452 -280 456 -170
rect 482 -280 486 -170
rect 452 -288 486 -280
rect 506 -170 540 -160
rect 506 -280 510 -170
rect 536 -280 540 -170
rect 856 -244 870 -240
rect 856 -254 860 -244
rect 864 -254 870 -244
rect 856 -258 870 -254
rect 886 -244 930 -240
rect 886 -254 900 -244
rect 916 -254 930 -244
rect 886 -258 930 -254
rect 946 -244 960 -240
rect 946 -254 952 -244
rect 956 -254 960 -244
rect 946 -258 960 -254
rect 1024 -244 1038 -240
rect 1024 -254 1028 -244
rect 1032 -254 1038 -244
rect 1024 -258 1038 -254
rect 1054 -244 1098 -240
rect 1054 -254 1068 -244
rect 1084 -254 1098 -244
rect 1054 -258 1098 -254
rect 1114 -244 1128 -240
rect 1114 -254 1120 -244
rect 1124 -254 1128 -244
rect 1114 -258 1128 -254
rect 506 -288 540 -280
<< pdiffusion >>
rect -48 474 -14 497
rect -48 120 -44 474
rect -21 120 -14 474
rect -48 113 -14 120
rect 6 474 40 497
rect 6 120 13 474
rect 36 120 40 474
rect 6 113 40 120
rect 856 504 870 518
rect 452 474 486 497
rect 452 120 456 474
rect 479 120 486 474
rect 452 113 486 120
rect 506 474 540 497
rect 506 120 513 474
rect 536 120 540 474
rect 506 113 540 120
rect 856 480 860 504
rect 866 480 870 504
rect 856 464 870 480
rect 886 510 930 518
rect 886 472 900 510
rect 916 472 930 510
rect 886 464 930 472
rect 946 504 960 518
rect 946 480 950 504
rect 956 480 960 504
rect 946 464 960 480
rect 1024 507 1038 522
rect 1024 483 1028 507
rect 1034 483 1038 507
rect 1024 468 1038 483
rect 1054 514 1098 522
rect 1054 476 1068 514
rect 1084 476 1098 514
rect 1054 468 1098 476
rect 1114 507 1128 522
rect 1114 483 1118 507
rect 1124 483 1128 507
rect 1114 468 1128 483
<< metal1 >>
rect 141 576 363 577
rect 641 576 825 577
rect 1140 576 1326 577
rect -157 556 1326 576
rect -118 502 -66 556
rect 58 502 110 556
rect 141 555 363 556
rect -66 120 -44 474
rect 13 106 36 120
rect 382 502 434 556
rect 558 502 610 556
rect 641 555 838 556
rect 882 555 934 556
rect 434 120 456 474
rect 513 106 536 120
rect 814 504 838 555
rect 838 480 860 504
rect 950 504 956 556
rect 1058 555 1110 556
rect 1140 551 1326 556
rect 1140 522 1158 551
rect 870 428 886 444
rect 900 405 916 472
rect 930 428 946 444
rect 1028 405 1034 483
rect 1038 436 1054 444
rect 1068 450 1084 476
rect 1098 436 1114 444
rect 1118 405 1124 483
rect 900 392 1124 405
rect -14 47 6 79
rect 14 47 36 106
rect 66 47 141 49
rect 486 47 506 79
rect 514 47 536 106
rect -122 27 6 47
rect -122 -40 -113 27
rect -14 -128 6 27
rect 10 46 141 47
rect 10 28 122 46
rect 137 28 141 46
rect 10 27 84 28
rect 408 27 506 47
rect 10 -170 36 27
rect 426 11 440 27
rect 486 -128 506 27
rect 510 42 809 47
rect 510 27 1062 42
rect 510 -170 536 27
rect 1268 23 1281 60
rect 808 -63 972 -62
rect 815 -72 972 -63
rect 870 -223 886 -208
rect 930 -223 946 -208
rect 952 -244 956 -206
rect 1038 -223 1054 -212
rect 1098 -223 1114 -213
rect 1120 -244 1124 -198
rect -44 -352 -18 -280
rect 456 -352 482 -280
rect 860 -330 864 -254
rect 1028 -322 1032 -254
rect 976 -330 1032 -322
rect 860 -340 1032 -330
rect 860 -352 982 -340
rect -44 -359 78 -352
rect -44 -422 -18 -359
rect 64 -422 78 -359
rect -44 -428 78 -422
rect -44 -444 -40 -428
rect -157 -458 -40 -444
rect -22 -458 56 -428
rect 74 -444 78 -428
rect 456 -359 578 -352
rect 860 -353 1078 -352
rect 456 -422 482 -359
rect 564 -422 578 -359
rect 456 -428 578 -422
rect 141 -444 363 -443
rect 456 -444 460 -428
rect 74 -458 460 -444
rect 478 -458 556 -428
rect 574 -444 578 -428
rect 956 -359 1078 -353
rect 956 -422 982 -359
rect 1064 -422 1078 -359
rect 956 -428 1078 -422
rect 956 -444 960 -428
rect 574 -458 960 -444
rect 978 -458 1056 -428
rect 1074 -444 1078 -428
rect 1074 -445 1148 -444
rect 1074 -458 1326 -445
rect -157 -463 1326 -458
rect -157 -464 648 -463
rect 843 -464 1326 -463
rect 141 -465 363 -464
rect 1136 -471 1326 -464
<< metal2 >>
rect 870 401 886 416
rect 870 394 874 401
rect 882 394 886 401
rect 870 392 886 394
rect 930 386 946 416
rect 930 380 934 386
rect 942 380 946 386
rect 930 377 946 380
rect 1038 382 1054 428
rect 1038 375 1042 382
rect 1050 375 1054 382
rect 1038 373 1054 375
rect 1068 82 1084 439
rect 1098 381 1114 428
rect 1098 375 1102 381
rect 1110 375 1114 381
rect 1098 372 1114 375
rect 952 76 1295 82
rect 952 60 1267 76
rect 1282 60 1295 76
rect 952 57 1295 60
rect 122 -17 137 28
rect 426 -10 440 1
rect 426 -15 430 -10
rect 436 -15 440 -10
rect 426 -17 440 -15
rect 122 -27 125 -17
rect 134 -27 137 -17
rect 122 -29 137 -27
rect 776 -28 906 -26
rect 776 -34 900 -28
rect 904 -34 906 -28
rect 776 -36 906 -34
rect -122 -96 -113 -48
rect 768 -64 808 -63
rect 777 -72 808 -64
rect 870 -180 886 -178
rect 870 -186 874 -180
rect 882 -186 886 -180
rect 870 -198 886 -186
rect 930 -180 946 -178
rect 930 -186 934 -180
rect 942 -186 946 -180
rect 930 -198 946 -186
rect 952 -198 956 57
rect 1073 38 1087 42
rect 1073 30 1080 38
rect 1084 30 1087 38
rect 1073 27 1087 30
rect 982 -65 1008 -62
rect 982 -69 999 -65
rect 1006 -69 1008 -65
rect 982 -72 1008 -69
rect 1038 -188 1043 -182
rect 1049 -188 1055 -182
rect 1038 -205 1055 -188
rect 1054 -212 1055 -205
rect 1098 -186 1103 -181
rect 1109 -186 1114 -181
rect 1098 -206 1114 -186
rect 1120 -189 1124 57
<< metal3 >>
rect 872 401 884 404
rect 872 394 874 401
rect 882 394 884 401
rect 427 -10 439 -6
rect 122 -17 137 -11
rect 122 -27 125 -17
rect 134 -27 137 -17
rect 122 -58 137 -27
rect 427 -15 430 -10
rect 436 -15 439 -10
rect 427 -21 439 -15
rect 427 -26 780 -21
rect 427 -36 768 -26
rect 776 -36 780 -26
rect 427 -39 780 -36
rect 122 -64 782 -58
rect 122 -72 768 -64
rect 777 -72 782 -64
rect 122 -76 782 -72
rect 872 -92 884 394
rect 932 386 944 390
rect 932 380 934 386
rect 942 380 944 386
rect 932 -26 944 380
rect 898 -28 944 -26
rect 898 -34 900 -28
rect 904 -34 944 -28
rect 898 -36 944 -34
rect -127 -96 884 -92
rect -127 -104 -122 -96
rect -113 -104 884 -96
rect -127 -108 884 -104
rect 872 -180 884 -108
rect 872 -186 874 -180
rect 882 -186 884 -180
rect 872 -188 884 -186
rect 932 -180 944 -36
rect 1040 382 1052 384
rect 1040 375 1042 382
rect 1050 375 1052 382
rect 1040 -62 1052 375
rect 1100 381 1112 384
rect 1100 375 1102 381
rect 1110 375 1112 381
rect 1100 40 1112 375
rect 1078 38 1112 40
rect 1078 30 1080 38
rect 1084 30 1112 38
rect 1078 28 1112 30
rect 996 -65 1052 -62
rect 996 -69 999 -65
rect 1006 -69 1052 -65
rect 996 -72 1052 -69
rect 932 -186 934 -180
rect 942 -186 944 -180
rect 932 -188 944 -186
rect 1040 -182 1052 -72
rect 1040 -188 1043 -182
rect 1049 -188 1052 -182
rect 1100 -181 1112 28
rect 1100 -186 1103 -181
rect 1109 -186 1112 -181
rect 1100 -188 1112 -186
rect 1040 -190 1052 -188
<< ntransistor >>
rect -14 -288 6 -160
rect 486 -288 506 -160
rect 870 -258 886 -240
rect 930 -258 946 -240
rect 1038 -258 1054 -240
rect 1098 -258 1114 -240
<< ptransistor >>
rect -14 113 6 497
rect 486 113 506 497
rect 870 464 886 518
rect 930 464 946 518
rect 1038 468 1054 522
rect 1098 468 1114 522
<< polycontact >>
rect -14 79 6 106
rect 870 444 886 452
rect 930 444 946 452
rect 1038 444 1054 452
rect 1098 444 1114 452
rect 486 79 506 106
rect -14 -152 6 -128
rect 486 -152 506 -128
rect 870 -234 886 -223
rect 930 -234 946 -223
rect 1038 -230 1054 -223
rect 1098 -230 1114 -223
<< ndcontact >>
rect -44 -280 -18 -170
rect 10 -280 36 -170
rect 456 -280 482 -170
rect 510 -280 536 -170
rect 860 -254 864 -244
rect 900 -254 916 -244
rect 952 -254 956 -244
rect 1028 -254 1032 -244
rect 1068 -254 1084 -244
rect 1120 -254 1124 -244
<< pdcontact >>
rect -44 120 -21 474
rect 13 120 36 474
rect 456 120 479 474
rect 513 120 536 474
rect 860 480 866 504
rect 900 472 916 510
rect 950 480 956 504
rect 1028 483 1034 507
rect 1068 476 1084 514
rect 1118 483 1124 507
<< m2contact >>
rect 870 416 886 428
rect 930 416 946 428
rect 1068 439 1084 450
rect 1038 428 1054 436
rect 1098 428 1114 436
rect 1267 60 1282 76
rect -122 -48 -113 -40
rect 122 28 137 46
rect 426 1 440 11
rect 1062 27 1073 42
rect 808 -72 815 -63
rect 972 -72 982 -62
rect 1120 -198 1124 -189
rect 870 -208 886 -198
rect 930 -208 946 -198
rect 952 -206 956 -198
rect 1038 -212 1054 -205
rect 1098 -213 1114 -206
<< m3contact >>
rect 874 394 882 401
rect 934 380 942 386
rect 1042 375 1050 382
rect 1102 375 1110 381
rect 430 -15 436 -10
rect 125 -27 134 -17
rect 768 -36 776 -26
rect 900 -34 904 -28
rect 768 -72 777 -64
rect -122 -104 -113 -96
rect 874 -186 882 -180
rect 934 -186 942 -180
rect 1080 30 1084 38
rect 999 -69 1006 -65
rect 1043 -188 1049 -182
rect 1103 -186 1109 -181
<< psubstratepcontact >>
rect -18 -422 64 -359
rect 482 -422 564 -359
rect 982 -422 1064 -359
rect -40 -458 -22 -428
rect 56 -458 74 -428
rect 460 -458 478 -428
rect 556 -458 574 -428
rect 960 -458 978 -428
rect 1056 -458 1074 -428
<< nsubstratencontact >>
rect -118 112 -66 502
rect 58 112 110 502
rect 382 112 434 502
rect 558 112 610 502
rect 814 480 838 504
rect 1140 472 1158 522
<< labels >>
rlabel metal1 -95 37 -95 37 1 B
rlabel metal1 424 36 424 36 1 A
rlabel metal1 334 565 334 565 1 Vdd
rlabel metal1 338 -456 338 -456 1 Gnd
rlabel metal1 1274 27 1274 27 1 Out
<< end >>
