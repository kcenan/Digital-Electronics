magic
tech scmos
timestamp 1494886329
<< nwell >>
rect -127 106 364 518
rect 432 106 677 518
rect 737 106 982 518
rect 1034 106 1525 518
rect 1585 106 2076 518
rect 2136 106 2381 518
rect 2441 106 2686 518
rect 2738 106 3229 518
<< polysilicon >>
rect -14 497 6 514
rect -14 106 6 113
rect 222 497 242 504
rect 222 400 242 407
rect 545 497 565 514
rect 545 106 565 113
rect 850 497 870 514
rect 850 106 870 113
rect 1147 497 1167 514
rect 1147 106 1167 113
rect 1383 497 1403 504
rect 1383 400 1403 407
rect 1698 497 1718 514
rect 1698 106 1718 113
rect 1934 497 1954 504
rect 1934 400 1954 407
rect 2249 497 2269 514
rect 2249 106 2269 113
rect 2554 497 2574 514
rect 2554 106 2574 113
rect 2851 497 2871 514
rect 2851 106 2871 113
rect 3087 497 3107 504
rect 3087 400 3107 407
rect -14 -160 6 -152
rect 545 -160 565 -152
rect 850 -160 870 -152
rect 1147 -160 1167 -152
rect 1698 -160 1718 -152
rect 2249 -160 2269 -152
rect 2554 -160 2574 -152
rect 2851 -160 2871 -152
rect -14 -299 6 -288
rect 222 -292 242 -282
rect 545 -299 565 -288
rect 850 -299 870 -288
rect 1147 -299 1167 -288
rect 1383 -292 1403 -282
rect 1698 -299 1718 -288
rect 1934 -292 1954 -282
rect 2249 -299 2269 -288
rect 2554 -299 2574 -288
rect 2851 -299 2871 -288
rect 3087 -292 3107 -282
rect 222 -327 242 -322
rect 1383 -327 1403 -322
rect 1934 -327 1954 -322
rect 3087 -327 3107 -322
<< ndiffusion >>
rect -48 -170 -14 -160
rect -48 -280 -44 -170
rect -18 -280 -14 -170
rect -48 -288 -14 -280
rect 6 -170 40 -160
rect 6 -280 10 -170
rect 36 -280 40 -170
rect 6 -288 40 -280
rect 511 -170 545 -160
rect 511 -280 515 -170
rect 541 -280 545 -170
rect 511 -288 545 -280
rect 565 -170 599 -160
rect 565 -280 569 -170
rect 595 -280 599 -170
rect 565 -288 599 -280
rect 816 -170 850 -160
rect 816 -280 820 -170
rect 846 -280 850 -170
rect 816 -288 850 -280
rect 870 -170 904 -160
rect 870 -280 874 -170
rect 900 -280 904 -170
rect 870 -288 904 -280
rect 1113 -170 1147 -160
rect 1113 -280 1117 -170
rect 1143 -280 1147 -170
rect 1113 -288 1147 -280
rect 1167 -170 1201 -160
rect 1167 -280 1171 -170
rect 1197 -280 1201 -170
rect 1167 -288 1201 -280
rect 1664 -170 1698 -160
rect 1664 -280 1668 -170
rect 1694 -280 1698 -170
rect 132 -296 222 -292
rect 132 -318 140 -296
rect 214 -318 222 -296
rect 132 -322 222 -318
rect 242 -296 330 -292
rect 242 -318 250 -296
rect 324 -318 330 -296
rect 1664 -288 1698 -280
rect 1718 -170 1752 -160
rect 1718 -280 1722 -170
rect 1748 -280 1752 -170
rect 1718 -288 1752 -280
rect 2215 -170 2249 -160
rect 2215 -280 2219 -170
rect 2245 -280 2249 -170
rect 1293 -296 1383 -292
rect 242 -322 330 -318
rect 1293 -318 1301 -296
rect 1375 -318 1383 -296
rect 1293 -322 1383 -318
rect 1403 -296 1491 -292
rect 1403 -318 1411 -296
rect 1485 -318 1491 -296
rect 2215 -288 2249 -280
rect 2269 -170 2303 -160
rect 2269 -280 2273 -170
rect 2299 -280 2303 -170
rect 2269 -288 2303 -280
rect 2520 -170 2554 -160
rect 2520 -280 2524 -170
rect 2550 -280 2554 -170
rect 2520 -288 2554 -280
rect 2574 -170 2608 -160
rect 2574 -280 2578 -170
rect 2604 -280 2608 -170
rect 2574 -288 2608 -280
rect 2817 -170 2851 -160
rect 2817 -280 2821 -170
rect 2847 -280 2851 -170
rect 2817 -288 2851 -280
rect 2871 -170 2905 -160
rect 2871 -280 2875 -170
rect 2901 -280 2905 -170
rect 2871 -288 2905 -280
rect 1844 -296 1934 -292
rect 1403 -322 1491 -318
rect 1844 -318 1852 -296
rect 1926 -318 1934 -296
rect 1844 -322 1934 -318
rect 1954 -296 2042 -292
rect 1954 -318 1962 -296
rect 2036 -318 2042 -296
rect 2997 -296 3087 -292
rect 1954 -322 2042 -318
rect 2997 -318 3005 -296
rect 3079 -318 3087 -296
rect 2997 -322 3087 -318
rect 3107 -296 3195 -292
rect 3107 -318 3115 -296
rect 3189 -318 3195 -296
rect 3107 -322 3195 -318
<< pdiffusion >>
rect -48 474 -14 497
rect -48 120 -44 474
rect -21 120 -14 474
rect -48 113 -14 120
rect 6 474 40 497
rect 6 120 13 474
rect 36 120 40 474
rect 6 113 40 120
rect 132 486 222 497
rect 132 416 140 486
rect 214 416 222 486
rect 132 407 222 416
rect 242 486 330 497
rect 242 416 250 486
rect 324 416 330 486
rect 242 407 330 416
rect 511 474 545 497
rect 511 120 515 474
rect 538 120 545 474
rect 511 113 545 120
rect 565 474 599 497
rect 565 120 572 474
rect 595 120 599 474
rect 565 113 599 120
rect 816 474 850 497
rect 816 120 820 474
rect 843 120 850 474
rect 816 113 850 120
rect 870 474 904 497
rect 870 120 877 474
rect 900 120 904 474
rect 870 113 904 120
rect 1113 474 1147 497
rect 1113 120 1117 474
rect 1140 120 1147 474
rect 1113 113 1147 120
rect 1167 474 1201 497
rect 1167 120 1174 474
rect 1197 120 1201 474
rect 1167 113 1201 120
rect 1293 486 1383 497
rect 1293 416 1301 486
rect 1375 416 1383 486
rect 1293 407 1383 416
rect 1403 486 1491 497
rect 1403 416 1411 486
rect 1485 416 1491 486
rect 1403 407 1491 416
rect 1664 474 1698 497
rect 1664 120 1668 474
rect 1691 120 1698 474
rect 1664 113 1698 120
rect 1718 474 1752 497
rect 1718 120 1725 474
rect 1748 120 1752 474
rect 1718 113 1752 120
rect 1844 486 1934 497
rect 1844 416 1852 486
rect 1926 416 1934 486
rect 1844 407 1934 416
rect 1954 486 2042 497
rect 1954 416 1962 486
rect 2036 416 2042 486
rect 1954 407 2042 416
rect 2215 474 2249 497
rect 2215 120 2219 474
rect 2242 120 2249 474
rect 2215 113 2249 120
rect 2269 474 2303 497
rect 2269 120 2276 474
rect 2299 120 2303 474
rect 2269 113 2303 120
rect 2520 474 2554 497
rect 2520 120 2524 474
rect 2547 120 2554 474
rect 2520 113 2554 120
rect 2574 474 2608 497
rect 2574 120 2581 474
rect 2604 120 2608 474
rect 2574 113 2608 120
rect 2817 474 2851 497
rect 2817 120 2821 474
rect 2844 120 2851 474
rect 2817 113 2851 120
rect 2871 474 2905 497
rect 2871 120 2878 474
rect 2901 120 2905 474
rect 2871 113 2905 120
rect 2997 486 3087 497
rect 2997 416 3005 486
rect 3079 416 3087 486
rect 2997 407 3087 416
rect 3107 486 3195 497
rect 3107 416 3115 486
rect 3189 416 3195 486
rect 3107 407 3195 416
<< metal1 >>
rect -157 556 3282 576
rect -118 502 -66 556
rect 58 502 110 556
rect 222 518 242 526
rect -66 120 -44 474
rect 13 106 36 120
rect 441 502 493 556
rect -14 74 6 79
rect -14 56 -12 74
rect -14 47 6 56
rect 14 47 36 106
rect -92 27 6 47
rect -92 -2 -80 16
rect -14 -128 6 27
rect 10 27 122 47
rect 10 -170 36 27
rect -44 -352 -18 -280
rect 106 -327 122 27
rect 140 16 214 416
rect 140 -2 158 16
rect 184 -2 214 16
rect 140 -296 214 -2
rect 250 16 324 416
rect 617 502 669 556
rect 493 120 515 474
rect 572 106 595 120
rect 746 502 798 556
rect 922 502 974 556
rect 798 120 820 474
rect 877 106 900 120
rect 1043 502 1095 556
rect 1219 502 1271 556
rect 1383 518 1403 526
rect 1095 120 1117 474
rect 1174 106 1197 120
rect 1594 502 1646 556
rect 545 47 565 79
rect 573 47 595 106
rect 850 47 870 79
rect 878 47 900 106
rect 1147 47 1167 79
rect 1175 47 1197 106
rect 467 27 565 47
rect 467 16 486 27
rect 250 -2 388 16
rect 414 -2 486 16
rect 250 -296 324 -2
rect 545 -128 565 27
rect 569 27 666 47
rect 688 27 870 47
rect 569 -170 595 27
rect 850 -128 870 27
rect 874 27 954 47
rect 1094 27 1167 47
rect 874 -170 900 27
rect 935 16 954 27
rect 935 -2 1081 16
rect 1147 -28 1167 27
rect 1147 -128 1167 -46
rect 1171 27 1227 47
rect 1171 -170 1197 27
rect 1301 16 1375 416
rect 1301 -2 1319 16
rect 1345 -2 1375 16
rect 106 -344 222 -327
rect 515 -352 541 -280
rect 820 -352 846 -280
rect 1117 -352 1143 -280
rect 1267 -327 1283 -46
rect 1301 -296 1375 -2
rect 1411 16 1485 416
rect 1770 502 1822 556
rect 1934 518 1954 526
rect 1646 120 1668 474
rect 1725 106 1748 120
rect 2145 502 2197 556
rect 1698 47 1718 79
rect 1726 47 1748 106
rect 1644 27 1718 47
rect 1411 -2 1516 16
rect 1411 -296 1485 -2
rect 1620 -62 1644 27
rect 1698 -28 1718 27
rect 1698 -128 1718 -46
rect 1722 27 1778 47
rect 1722 -170 1748 27
rect 1852 16 1926 416
rect 1852 -2 1870 16
rect 1896 -2 1926 16
rect 1267 -344 1383 -327
rect 1668 -352 1694 -280
rect 1818 -327 1834 -46
rect 1852 -296 1926 -2
rect 1962 16 2036 416
rect 2321 502 2373 556
rect 2197 120 2219 474
rect 2276 106 2299 120
rect 2450 502 2502 556
rect 2626 502 2678 556
rect 2502 120 2524 474
rect 2581 106 2604 120
rect 2747 502 2799 556
rect 2923 502 2975 556
rect 3087 518 3107 526
rect 2799 120 2821 474
rect 2878 106 2901 120
rect 2249 47 2269 79
rect 2277 47 2299 106
rect 2554 47 2574 79
rect 2582 47 2604 106
rect 2851 72 2871 79
rect 2851 47 2871 55
rect 2879 47 2901 106
rect 2171 27 2269 47
rect 2171 16 2190 27
rect 1962 -2 2082 16
rect 2106 -2 2190 16
rect 1962 -296 2036 -2
rect 2249 -128 2269 27
rect 2273 27 2574 47
rect 2273 -170 2299 27
rect 2554 -32 2574 27
rect 2554 -128 2574 -54
rect 2578 27 2710 47
rect 2795 27 2871 47
rect 2578 -170 2604 27
rect 2690 16 2710 27
rect 2690 -2 2785 16
rect 2851 -128 2871 27
rect 2875 27 2987 47
rect 2875 -170 2901 27
rect 1818 -344 1934 -327
rect 2219 -352 2245 -280
rect 2524 -352 2550 -280
rect 2821 -352 2847 -280
rect 2971 -327 2987 27
rect 3005 16 3079 416
rect 3005 -2 3023 16
rect 3049 -2 3079 16
rect 3005 -296 3079 -2
rect 3115 16 3189 416
rect 3230 38 3252 60
rect 3115 -2 3210 16
rect 3115 -296 3189 -2
rect 2971 -344 3087 -327
rect -44 -357 198 -352
rect -44 -422 -31 -357
rect 189 -422 198 -357
rect -44 -428 198 -422
rect -44 -444 -40 -428
rect -157 -458 -40 -444
rect -22 -458 56 -428
rect 74 -444 198 -428
rect 515 -359 637 -352
rect 515 -422 541 -359
rect 623 -422 637 -359
rect 515 -428 637 -422
rect 515 -444 519 -428
rect 74 -458 519 -444
rect 537 -458 615 -428
rect 633 -444 637 -428
rect 820 -359 942 -352
rect 820 -422 846 -359
rect 928 -422 942 -359
rect 820 -428 942 -422
rect 820 -444 824 -428
rect 633 -458 824 -444
rect 842 -458 920 -428
rect 938 -444 942 -428
rect 1117 -357 1359 -352
rect 1117 -422 1130 -357
rect 1350 -422 1359 -357
rect 1117 -428 1359 -422
rect 1117 -444 1121 -428
rect 938 -458 1121 -444
rect 1139 -458 1217 -428
rect 1235 -444 1359 -428
rect 1668 -357 1910 -352
rect 1668 -422 1681 -357
rect 1901 -422 1910 -357
rect 1668 -428 1910 -422
rect 1668 -444 1672 -428
rect 1235 -458 1672 -444
rect 1690 -458 1768 -428
rect 1786 -444 1910 -428
rect 2219 -359 2341 -352
rect 2219 -422 2245 -359
rect 2327 -422 2341 -359
rect 2219 -428 2341 -422
rect 2219 -444 2223 -428
rect 1786 -458 2223 -444
rect 2241 -458 2319 -428
rect 2337 -444 2341 -428
rect 2524 -359 2646 -352
rect 2524 -422 2550 -359
rect 2632 -422 2646 -359
rect 2524 -428 2646 -422
rect 2524 -444 2528 -428
rect 2337 -458 2528 -444
rect 2546 -458 2624 -428
rect 2642 -444 2646 -428
rect 2821 -357 3063 -352
rect 2821 -422 2834 -357
rect 3054 -422 3063 -357
rect 2821 -428 3063 -422
rect 2821 -444 2825 -428
rect 2642 -458 2825 -444
rect 2843 -458 2921 -428
rect 2939 -444 3063 -428
rect 2939 -458 3282 -444
rect -157 -464 3282 -458
<< metal2 >>
rect 66 526 222 542
rect 1227 526 1383 542
rect 1778 526 1934 542
rect 2931 526 3087 542
rect 66 74 84 526
rect 6 56 1010 74
rect 1034 56 1094 74
rect -66 -2 158 16
rect 388 -94 414 -2
rect 666 -62 688 27
rect 1010 -6 1034 56
rect 1069 47 1094 56
rect 1227 47 1245 526
rect 1448 58 1644 78
rect 1095 -2 1319 16
rect 1448 -6 1470 58
rect 1620 47 1644 58
rect 1010 -24 1470 -6
rect 1478 26 1580 44
rect 1778 47 1796 526
rect 2931 72 2949 526
rect 2871 55 2949 72
rect 1940 27 2773 47
rect 3084 38 3211 60
rect 1167 -46 1267 -28
rect 1478 -62 1500 26
rect 1560 16 1580 26
rect 666 -84 1500 -62
rect 1560 -2 1870 16
rect 1516 -94 1538 -2
rect 1718 -46 1818 -28
rect 1940 -62 1964 27
rect 1662 -84 1964 -62
rect 2799 -2 3023 16
rect 388 -116 1538 -94
rect 2082 -96 2106 -2
rect 3084 -32 3110 38
rect 2574 -54 3110 -32
rect 3210 -96 3232 -2
rect 2082 -117 3232 -96
<< ntransistor >>
rect -14 -288 6 -160
rect 545 -288 565 -160
rect 850 -288 870 -160
rect 1147 -288 1167 -160
rect 222 -322 242 -292
rect 1698 -288 1718 -160
rect 1383 -322 1403 -292
rect 2249 -288 2269 -160
rect 2554 -288 2574 -160
rect 2851 -288 2871 -160
rect 1934 -322 1954 -292
rect 3087 -322 3107 -292
<< ptransistor >>
rect -14 113 6 497
rect 222 407 242 497
rect 545 113 565 497
rect 850 113 870 497
rect 1147 113 1167 497
rect 1383 407 1403 497
rect 1698 113 1718 497
rect 1934 407 1954 497
rect 2249 113 2269 497
rect 2554 113 2574 497
rect 2851 113 2871 497
rect 3087 407 3107 497
<< polycontact >>
rect 222 504 242 518
rect -14 79 6 106
rect 545 79 565 106
rect 1383 504 1403 518
rect 850 79 870 106
rect 1934 504 1954 518
rect 1147 79 1167 106
rect 1698 79 1718 106
rect 2249 79 2269 106
rect 3087 504 3107 518
rect 2554 79 2574 106
rect 2851 79 2871 106
rect -14 -152 6 -128
rect 545 -152 565 -128
rect 850 -152 870 -128
rect 1147 -152 1167 -128
rect 1698 -152 1718 -128
rect 2249 -152 2269 -128
rect 2554 -152 2574 -128
rect 2851 -152 2871 -128
rect 222 -344 242 -327
rect 1383 -344 1403 -327
rect 1934 -344 1954 -327
rect 3087 -344 3107 -327
<< ndcontact >>
rect -44 -280 -18 -170
rect 10 -280 36 -170
rect 515 -280 541 -170
rect 569 -280 595 -170
rect 820 -280 846 -170
rect 874 -280 900 -170
rect 1117 -280 1143 -170
rect 1171 -280 1197 -170
rect 1668 -280 1694 -170
rect 140 -318 214 -296
rect 250 -318 324 -296
rect 1722 -280 1748 -170
rect 2219 -280 2245 -170
rect 1301 -318 1375 -296
rect 1411 -318 1485 -296
rect 2273 -280 2299 -170
rect 2524 -280 2550 -170
rect 2578 -280 2604 -170
rect 2821 -280 2847 -170
rect 2875 -280 2901 -170
rect 1852 -318 1926 -296
rect 1962 -318 2036 -296
rect 3005 -318 3079 -296
rect 3115 -318 3189 -296
<< pdcontact >>
rect -44 120 -21 474
rect 13 120 36 474
rect 140 416 214 486
rect 250 416 324 486
rect 515 120 538 474
rect 572 120 595 474
rect 820 120 843 474
rect 877 120 900 474
rect 1117 120 1140 474
rect 1174 120 1197 474
rect 1301 416 1375 486
rect 1411 416 1485 486
rect 1668 120 1691 474
rect 1725 120 1748 474
rect 1852 416 1926 486
rect 1962 416 2036 486
rect 2219 120 2242 474
rect 2276 120 2299 474
rect 2524 120 2547 474
rect 2581 120 2604 474
rect 2821 120 2844 474
rect 2878 120 2901 474
rect 3005 416 3079 486
rect 3115 416 3189 486
<< m2contact >>
rect 222 526 242 542
rect -12 56 6 74
rect -80 -2 -66 16
rect 158 -2 184 16
rect 1383 526 1403 542
rect 1010 56 1034 74
rect 388 -2 414 16
rect 666 27 688 47
rect 1069 27 1094 47
rect 1081 -2 1095 16
rect 1147 -46 1167 -28
rect 1227 27 1245 47
rect 1319 -2 1345 16
rect 1267 -46 1283 -28
rect 1934 526 1954 542
rect 1620 27 1644 47
rect 1516 -2 1538 16
rect 1698 -46 1718 -28
rect 1620 -84 1662 -62
rect 1778 27 1796 47
rect 1870 -2 1896 16
rect 1818 -46 1834 -28
rect 3087 526 3107 542
rect 2851 55 2871 72
rect 2082 -2 2106 16
rect 2554 -54 2574 -32
rect 2773 27 2795 47
rect 2785 -2 2799 16
rect 3023 -2 3049 16
rect 3211 38 3230 60
rect 3210 -2 3232 16
<< psubstratepcontact >>
rect -31 -422 189 -357
rect 541 -422 623 -359
rect 846 -422 928 -359
rect 1130 -422 1350 -357
rect 1681 -422 1901 -357
rect 2245 -422 2327 -359
rect 2550 -422 2632 -359
rect 2834 -422 3054 -357
rect -40 -458 -22 -428
rect 56 -458 74 -428
rect 519 -458 537 -428
rect 615 -458 633 -428
rect 824 -458 842 -428
rect 920 -458 938 -428
rect 1121 -458 1139 -428
rect 1217 -458 1235 -428
rect 1672 -458 1690 -428
rect 1768 -458 1786 -428
rect 2223 -458 2241 -428
rect 2319 -458 2337 -428
rect 2528 -458 2546 -428
rect 2624 -458 2642 -428
rect 2825 -458 2843 -428
rect 2921 -458 2939 -428
<< nsubstratencontact >>
rect -118 112 -66 502
rect 58 112 110 502
rect 441 112 493 502
rect 617 112 669 502
rect 746 112 798 502
rect 922 112 974 502
rect 1043 112 1095 502
rect 1219 112 1271 502
rect 1594 112 1646 502
rect 1770 112 1822 502
rect 2145 112 2197 502
rect 2321 112 2373 502
rect 2450 112 2502 502
rect 2626 112 2678 502
rect 2747 112 2799 502
rect 2923 112 2975 502
<< labels >>
rlabel metal1 1156 566 1156 566 1 vdd!
rlabel metal1 1157 -454 1157 -454 1 gnd!
rlabel metal1 -88 37 -88 37 1 clk
rlabel metal1 3245 50 3245 50 1 out
rlabel metal1 -87 7 -87 7 1 in
<< end >>
