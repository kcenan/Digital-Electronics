* SPICE3 file created from inv4x.ext - technology: scmos

m1000 out in vdd vdd pfet w=96u l=20u
+ ad=3264p pd=260u as=3264p ps=260u 
m1001 out in gnd Gnd nfet w=32u l=20u
+ ad=1088p pd=132u as=1088p ps=132u 
C0 vdd in 46.4fF
C1 vdd out 42.2fF
C2 gnd GND 464.4fF
C3 out GND 464.4fF
C4 in GND 438.2fF
C5 vdd GND 1414.5fF
